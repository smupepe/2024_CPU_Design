module pipeline(

);



endmodule